/*
 -- ============================================================================
 -- FILE NAME	: nettype.h
 -- DESCRIPTION : デフォルトネットタイプの指定
 -- ----------------------------------------------------------------------------
 -- Revision  Date		  Coding_by	 Comment
 -- 1.0.0	  2011/04/26  suito		 新規作成
 -- ============================================================================
*/

`ifndef __NETTYPE_HEADER__	   // インクルードガード
	`define __NETTYPE_HEADER__

	/********** デフォルトネットタイプ : いずれか1つを選択 **********/
	`default_nettype none	   // none (推奨)
//	`default_nettype wire	   // wire (Verilog標準)

`endif
